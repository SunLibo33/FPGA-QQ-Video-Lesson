library verilog;
use verilog.vl_types.all;
entity tb_ex_spi is
end tb_ex_spi;
