library verilog;
use verilog.vl_types.all;
entity tb_ex_fsm is
end tb_ex_fsm;
