library verilog;
use verilog.vl_types.all;
entity tb_ex_case is
end tb_ex_case;
