`timescale 1ns/100ps

module tb_ex_fifo();

reg tb_w_clk;  
reg tb_r_clk;  
reg tb_rst_n;  
reg tb_w_en;   
reg [7:0]tb_w_data;
reg tb_r_en;
 
wire tb_w_full;   
wire [7:0]tb_r_data; 
wire tb_r_empty;

parameter CLK_P=20;

initial
  begin
  	tb_w_clk=1'b0;
  	tb_r_clk=1'b0;
  	tb_rst_n=1'b0;
  	#200
  	tb_rst_n=1'b1;
  end
 
initial
  begin
  	tb_w_en=1'b0;
  	tb_w_data=8'h00;
    #300
    write_data(258);
  end  

initial
  begin
  	tb_r_en=1'b0;
  	@(posedge tb_w_full)
  	#40;
  	read_data(256);
 
  end   
  
always #(CLK_P/2) tb_w_clk=~tb_w_clk;
always #(CLK_P/2) tb_r_clk=~tb_r_clk;

ex_fifo ex_fifo_instance(
       .w_clk  (tb_w_clk  ) ,
       .r_clk  (tb_r_clk  ) ,
       .rst_n  (tb_rst_n  ) ,
       .w_en   (tb_w_en   ) ,
       .w_data (tb_w_data ) ,
       .w_full (tb_w_full ) ,
       .r_en   (tb_r_en   ) ,
       .r_data (tb_r_data ) ,
       .r_empty(tb_r_empty)
);


task write_data(len);
     integer i,len;
     begin
     	 for(i=0;i<len;i=i+1)
     	   begin
     	   	@(posedge tb_w_clk);
     	   	   tb_w_en=1'b1;
  	         tb_w_data=i;
     	   end
     	 @(posedge tb_w_clk);
  	     tb_w_en=1'b0;
  	     tb_w_data=8'h00;     	 
     end

endtask

task read_data(len);
     integer i,len;
     begin
     	 for(i=0;i<len;i=i+1)
     	   begin
     	   	@(posedge tb_r_clk);
     	   	   tb_r_en=1'b1;
     	   end
     	 @(posedge tb_w_clk);
  	     tb_r_en=1'b0;    	 
     end

endtask

endmodule
   