library verilog;
use verilog.vl_types.all;
entity TB_SPI is
end TB_SPI;
