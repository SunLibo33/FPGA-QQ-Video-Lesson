library verilog;
use verilog.vl_types.all;
entity tb_ex_shift_reg is
end tb_ex_shift_reg;
